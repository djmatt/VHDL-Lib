--------------------------------------------------------------------------------------------------
--        FIR Filter Testbench
--------------------------------------------------------------------------------------------------
-- Matthew Dallmeyer - d01matt@gmail.com

--------------------------------------------------------------------------------------------------
--        ENTITY
--------------------------------------------------------------------------------------------------
library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;

library work;
   use work.tb_clockgen_pkg.all;
   use work.tb_read_csv_pkg.all;
   use work.tb_write_csv_pkg.all;
   use work.dsp_pkg.all;
   use work.sparse_fir_filter_pkg.all;

--This module is a test-bench for simulating the fir filter
entity tb_sparse_fir_filter is
end tb_sparse_fir_filter;

--------------------------------------------------------------------------------------------------
--        ARCHITECTURE
--------------------------------------------------------------------------------------------------
architecture sim of tb_sparse_fir_filter is

   constant INPUT_FILE  : string 
      := "X:\Education\Masters Thesis\matlab\sparse_fir_filter\chirp.csv";
   
--   constant TEST_FILTER : coefficient_array  := LOW_PASS_21;
--   constant OUTPUT_FILE : string 
--      := "X:\Education\Masters Thesis\matlab\sparse_fir_filter\chirp_lowpass21.csv";  
   
--   constant TEST_FILTER : coefficient_array  := HIGH_PASS_41;
--   constant OUTPUT_FILE : string 
--      := "X:\Education\Masters Thesis\matlab\sparse_fir_filter\chirp_highpass41.csv";  
   
   constant TEST_FILTER : coefficient_array  := LOW_PASS_101;
   constant OUTPUT_FILE : string 
      := "X:\Education\Masters Thesis\matlab\sparse_fir_filter\chirp_lowpass101.csv";  
  
   signal rst        : std_logic := '0';
   signal clk        : std_logic := '0';
   signal sig        : std_logic_vector(NUM_SIG_BITS-1 downto 0) := (others => '0');
   signal filtered   : fir_sig := (others => '0');
begin

   --Instantiate clock generator
   clk1 : tb_clockgen
      generic map(PERIOD      => 10ns,
                  DUTY_CYCLE  => 0.50)
      port map(   clk         => clk);
      
   
   --Instantiate file reader
   reader : tb_read_csv
      generic map(FILENAME => INPUT_FILE)
      port map(   clk      => clk,
                  data     => sig);
   

   --Instantiate unit under test
   uut : entity work.sparse_fir_filter(behave)
      generic map(h    => TEST_FILTER)
      port map(   clk  => clk,
                  rst  => rst,
                  x    => signed(sig),
                  y    => filtered);
                                    
   --Instantiate a file writer
   writer : tb_write_csv
      generic map(FILENAME => OUTPUT_FILE)
      port map(   clk      => clk,
                  data     => std_logic_vector(filtered(30 downto 15)));

   --Main Process
   --TODO: Add a check for end of file, once reached terminate simulation.
   main: process
   begin
      rst <= '1';
      wait for 10ns;
      rst <= '0';
      wait;
   end process;
end sim;
