----------------------------------------------------------------------------------------------------
--        Digital Signal Processing package
----------------------------------------------------------------------------------------------------
-- Matthew Dallmeyer - d01matt@gmail.com

----------------------------------------------------------------------------------------------------
--        PACKAGE
----------------------------------------------------------------------------------------------------
library ieee;
   use ieee.std_logic_1164.all;
   use ieee.numeric_std.all;

package dsp_pkg is
   --Definitions for coefficients
   constant NUM_COEF_BITS : positive := 16;
   subtype coefficient is signed(NUM_COEF_BITS-1 downto 0);
   type coefficient_array is array (natural range <>) of coefficient;

   --Definitions for signal data
   constant NUM_SIG_BITS : positive := 16;
   subtype sig is signed(NUM_SIG_BITS-1 downto 0);
   subtype summed_sig is signed(NUM_SIG_BITS downto 0); --for when 2 sigs are added together
   constant NUM_SUMMED_SIG_BITS : positive := NUM_SIG_BITS+1;
   type sig_array is array (natural range <>) of sig;
   
   --Types for fir signal data - for use for internal FIR calculations
   --The size is based on the number of bits needed for calculation.  The multiplication of 
   --coefficient and signal is 16-bits + 16-bits.  The cumulative addtion of N taps will need 
   --require a log2(N) addtional bits.  Allowing for up to 256 taps, the full size will be 
   --16 + 16 + log2(256) or 40 bits
   constant MAX_TAPS : positive := 256;
   constant NUM_ADDED_TAPS_BITS : positive := 8; --log2(256)
   constant NUM_FIR_BITS : positive := NUM_COEF_BITS + NUM_SIG_BITS + NUM_ADDED_TAPS_BITS;
   subtype fir_sig is signed(NUM_FIR_BITS-1 downto 0);
   type fir_sig_array is array (natural range <>) of fir_sig;
   
   --Coefficients for FIR filters
   constant ZERO_COEF   : coefficient       := x"0000";
   
   constant LOW_PASS    : coefficient_array := (x"0000",
                                                x"0070",
                                                x"0000",
                                                x"fe7b",
                                                x"0000",
                                                x"0453",
                                                x"0000",
                                                x"f512",
                                                x"0000",
                                                x"27c2",
                                                x"4010",
                                                x"27c2",
                                                x"0000",
                                                x"f512",
                                                x"0000",
                                                x"0453",
                                                x"0000",
                                                x"fe7b",
                                                x"0000",
                                                x"0070",
                                                x"0000");
                                                
   constant HIGH_PASS   : coefficient_array := (x"0000",
                                                x"ff90",
                                                x"0000",
                                                x"0185",
                                                x"0000",
                                                x"fbad",
                                                x"0000",
                                                x"0aee",
                                                x"0000",
                                                x"d83e",
                                                x"4010",
                                                x"d83e",
                                                x"0000",
                                                x"0aee",
                                                x"0000",
                                                x"fbad",
                                                x"0000",
                                                x"0185",
                                                x"0000",
                                                x"ff90",
                                                x"0000");
                                                                                                
   constant PASS_THRU   : coefficient_array := (x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"3FFF",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000",
                                                x"0000");
   
   --Function declarations
--   type slice_type is array(natural range <>) of integer;
   function slice_coefficient_array (  original_array : coefficient_array; 
                                       num_cuts       : integer;
                                       cut            : integer) return coefficient_array;
   
end package;
 
----------------------------------------------------------------------------------------------------
--        PACKAGE BODY
----------------------------------------------------------------------------------------------------
library ieee;
   use ieee.std_logic_1164.all;

   
package body dsp_pkg is
   
   --This function slices a coefficient array into the polyphase slice of that array.
   --The original array is the coefficient array to be sliced
   --num_cuts is the number of sub-arrays that can be created
   --cut is the 1-based identifier of the cut desired (e.g. when num_cuts is 2, cut can be 1 or 2)
   function slice_coefficient_array (  original_array : coefficient_array; 
                                       num_cuts       : integer;
                                       cut            : integer) return coefficient_array is
      
      constant slice_len   : integer := (original_array'length - cut-1 + num_cuts) / num_cuts;
      constant result_len  : integer := (original_array'length - 1 + num_cuts) / num_cuts;
      variable result      : coefficient_array(1 to result_len)  := (others => (others => '0'));
   begin
      for index in 1 to slice_len loop
         result(index) := original_array(cut-1 + ((index-1)*num_cuts));
      end loop;
      return result;
   end function;
   
end package body;